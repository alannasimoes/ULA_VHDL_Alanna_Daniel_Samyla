LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY OPERACAO_DESLOCAR4BITS_ESQUERDA IS
    PORT (
        A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END OPERACAO_DESLOCAR4BITS_ESQUERDA;

ARCHITECTURE BEHAVIORAL OF OPERACAO_DESLOCAR4BITS_ESQUERDA IS
BEGIN
    PROCESS(A)
    BEGIN
        -- DESLOCAMENTO � ESQUERDA
        Z <= A(2 DOWNTO 0) & '0';
    END PROCESS;
END BEHAVIORAL;
