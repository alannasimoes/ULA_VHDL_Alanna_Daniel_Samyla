--------------------------------------------------------------------------------
-- COMPANY: 
-- ENGINEER:
--
-- CREATE DATE:   18:13:59 05/31/2024
-- DESIGN NAME:   
-- MODULE NAME:   C:/USERS/DANIEL/DESKTOP/SD/ULA_FINAL/TB_OPERACAO_SUBTRATOR4BITS.VHD
-- PROJECT NAME:  ULA_FINAL
-- TARGET DEVICE:  
-- TOOL VERSIONS:  
-- DESCRIPTION:   
-- 
-- VHDL TEST BENCH CREATED BY ISE FOR MODULE: OPERACAO_SUBTRATOR4BITS
-- 
-- DEPENDENCIES:
-- 
-- REVISION:
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS:
--
-- NOTES: 
-- THIS TESTBENCH HAS BEEN AUTOMATICALLY GENERATED USING TYPES STD_LOGIC AND
-- STD_LOGIC_VECTOR FOR THE PORTS OF THE UNIT UNDER TEST.  XILINX RECOMMENDS
-- THAT THESE TYPES ALWAYS BE USED FOR THE TOP-LEVEL I/O OF A DESIGN IN ORDER
-- TO GUARANTEE THAT THE TESTBENCH WILL BIND CORRECTLY TO THE POST-IMPLEMENTATION 
-- SIMULATION MODEL.
--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 
-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;
 
ENTITY TB_OPERACAO_SUBTRATOR4BITS IS
END TB_OPERACAO_SUBTRATOR4BITS;
 
ARCHITECTURE BEHAVIOR OF TB_OPERACAO_SUBTRATOR4BITS IS 
 
    -- COMPONENT DECLARATION FOR THE UNIT UNDER TEST (UUT)
 
    COMPONENT OPERACAO_SUBTRATOR4BITS
    PORT(
         A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         B : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         Z : OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
         CARRY_OUT : OUT  STD_LOGIC
        );
    END COMPONENT;
    

   --INPUTS
   SIGNAL A : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
   SIGNAL B : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');

 	--OUTPUTS
   SIGNAL Z : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL CARRY_OUT : STD_LOGIC;
   -- NO CLOCKS DETECTED IN PORT LIST. REPLACE <CLOCK> BELOW WITH 
   -- APPROPRIATE PORT NAME 
 
BEGIN
 
	-- INSTANTIATE THE UNIT UNDER TEST (UUT)
   UUT: OPERACAO_SUBTRATOR4BITS PORT MAP (
          A => A,
          B => B,
          Z => Z,
          CARRY_OUT => CARRY_OUT
        );

   -- STIMULUS PROCESS
   STIM_PROC: PROCESS
   BEGIN
		A <= "0100";
		B <= "0010";
      WAIT FOR 100 NS;
		A <= "0101";
		B <= "0011";
		WAIT FOR 100 NS;
		A <= "1111";
		B <= "1111";
   END PROCESS;

END;
