LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------------------------------
-------------------------------------ENTIDADE--------------------------------------
-----------------------------------------------------------------------------------
ENTITY ULA IS
    PORT (
        A_ULA : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        B_ULA : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        SEL_ULA : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        RESULTADO_ULA : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		  FLAG_CARRY_OUT_ULA : OUT STD_LOGIC;
		  FLAG_RESULTADO_NULO_ULA : OUT STD_LOGIC;
		  FLAG_OVERFLOW_ULA : OUT STD_LOGIC;
		  FLAG_RESULTADO_NEGATIVO_ULA : OUT  STD_LOGIC
    );
END ULA;
-------------------------------------------------------------------------------
----------------------------------ARQUITETURA----------------------------------
-------------------------------------------------------------------------------
ARCHITECTURE BEHAVIORAL OF ULA IS


--- IMPORTAR COMPONENTES PARA DENTRO DA ULA PARA PODER US-LOS NAS OPERAES
-------------------------------------------------------------------------------
---------------------------DECLARACAO DE COMPONENTES---------------------------
-------------------------------------------------------------------------------
COMPONENT MUX_8ENTRADAS IS
PORT(
        INPUT_0 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_1 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_2 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_3 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_4 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_5 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_6 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        INPUT_7 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        SEL     : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        OUTPUT  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END COMPONENT;

COMPONENT OPERACAO_AND IS
			PORT(
			A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT OPERACAO_OR IS
			PORT(
			A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT OPERACAO_XOR IS
			PORT(
			A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT OPERACAO_NOT IS
			PORT(
			A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT OPERACAO_SOMAR4BITS IS
	PORT(
        A, B        : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        CARRY_IN    : IN  STD_LOGIC;
        Z           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        CARRY_OUT   : OUT STD_LOGIC;
		  FLAG_RESULTADO_NULO : OUT STD_LOGIC;
        FLAG_OVERFLOW       : OUT STD_LOGIC);
END COMPONENT;

COMPONENT OPERACAO_SUBTRAIR4BITS IS
    PORT (
        A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        B : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        CARRY_OUT : OUT STD_LOGIC;
		  FLAG_RESULTADO_NEGATIVO : OUT STD_LOGIC);
END COMPONENT;

COMPONENT OPERACAO_DESLOCAR4BITS_ESQUERDA IS
    PORT (
        A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT OPERACAO_COMPARADOR_4BITS IS
    PORT (
        A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        B : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)); 
END COMPONENT;
 
---------------------------------------------------------------
---------------------SINAIS INTERMEDIARIOS---------------------
---------------------------------------------------------------
SIGNAL RESULTADO_OPERACAO : STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL RESULTADO_AND, 
RESULTADO_OR, 
RESULTADO_NOT, 
RESULTADO_XOR,
RESULTADO_SOMA,
RESULTADO_SUBTRACAO,
RESULTADO_COMPARADOR,
RESULTADO_DESLOCADOR: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

---------------------------------------------------------------
--------------------------INSTANCIAS---------------------------
---------------------------------------------------------------

--- AQUI EU ESTOU FAZENDO O PORT MAP DOS COMPONENTES PARA PODER USA-LOS NA ULA
--- BASICAMENTE A IDEIA  REUTILIZAR OS COMPONENTES, CRIAR SINAIS INTERMEDIARIOS E ENVIA-LOS AO MULTIPLEXADOR


--            		 							 _________________________
--           									|                         |
---RESULTADO_AND---(INPUT_0)-----------|                         |
---RESULTADO_OR---(INPUT_1)------------|                         |
---RESULTADO_NOT---(INPUT_2)-----------|                         |
---RESULTADO_XOR---(INPUT_3)-----------|       MULTIPLEXADOR     |
---RESULTADO_SOMA---(INPUT_4)----------|         8 PARA 1        |------(OUTPUT)------>(RESULTADO_ULA)
---RESULTADO_SUBTRACAO---(INPUT_5)-----|                         |
---RESULTADO_COMPARADOR---(INPUT_6)----|                         |
---RESULTADO_DESLOCADOR---(INPUT_7)----|_________________________|
							
														 --(SEL) = SEL_ULA


--- INSTANCIA DO COMPONENTE AND
      INSTANCIA_AND : OPERACAO_AND 
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					Z => RESULTADO_AND);
		
--- INSTANCIA DO COMPONENTE OR
      INSTANCIA_OR : OPERACAO_OR 
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					Z => RESULTADO_OR);

--- INSTANCIA DO COMPONENTE NOT
      INSTANCIA_NOT : OPERACAO_NOT
		PORT MAP (
					A => A_ULA,
					Z => RESULTADO_NOT);

					
--- INSTANCIA DO COMPONENTE XOR
      INSTANCIA_XOR : OPERACAO_XOR
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					Z => RESULTADO_XOR);

--- INSTANCIA DO COMPONENTE SOMADOR
      INSTANCIA_SOMADOR : OPERACAO_SOMAR4BITS 
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					CARRY_IN => '0',
					CARRY_OUT => FLAG_CARRY_OUT_ULA,
					Z => RESULTADO_SOMA,
					FLAG_RESULTADO_NULO => FLAG_RESULTADO_NULO_ULA,
					FLAG_OVERFLOW       => FLAG_OVERFLOW_ULA);

--- INSTANCIA DO COMPONENTE SUBTRATOR
      INSTANCIA_SUBTRATOR : OPERACAO_SUBTRAIR4BITS
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					CARRY_OUT => OPEN,
					Z => RESULTADO_SUBTRACAO,
					FLAG_RESULTADO_NEGATIVO => FLAG_RESULTADO_NEGATIVO_ULA);

--- INSTANCIA DO COMPONENTE COMPARADOR
      INSTANCIA_COMPARADOR : OPERACAO_COMPARADOR_4BITS
		PORT MAP (
					A => A_ULA,
					B => B_ULA,
					Z => RESULTADO_COMPARADOR);
					
--- INSTANCIA DO COMPONENTE DESLOCADOR (DESLOCA 1 BIT APESAR DO NOME)
      INSTANCIA_DESLOCADOR : OPERACAO_DESLOCAR4BITS_ESQUERDA
		PORT MAP (
					A => A_ULA,
					Z => RESULTADO_DESLOCADOR);
					
--- INSTANCIA DO MULTIPLEXADOR
		INSTANCIA_MULTIPLEXADOR : MUX_8ENTRADAS
		PORT MAP (
		  INPUT_0 => RESULTADO_AND,					--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO AND --> SEL_ULA = 000
        INPUT_1 => RESULTADO_OR,						--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO OR --> SELECT 001
        INPUT_2 => RESULTADO_NOT,					--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO NOT --> SELECT 010
        INPUT_3 => RESULTADO_XOR,					--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO XOR --> SELECT 011
        INPUT_4 => RESULTADO_SOMA,					--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO SOMA --> SELECT 100
        INPUT_5 => RESULTADO_SUBTRACAO,			--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO SUBTRACAO --> SELECT 101
        INPUT_6 => RESULTADO_COMPARADOR,			--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO COMPARACAO --> SELECT 110
        INPUT_7 => RESULTADO_DESLOCADOR,			--- SINAL INTERMEDIARIO QUE REPRESENTA O RESULTADO DA OPERACAO DESLOCAMENTO --> SELECT 111
        SEL     => SEL_ULA,							--- SINAL INTERMEDIARIO QUE REPRESENTA NOSSA ESCOLHA DE SAIDA DO MULTIPLEXADOR
        OUTPUT  => RESULTADO_ULA);					--- SINAL INTERMEDIARIO QUE REPRESENTA QUAL OPERACAO VAI SAIR NA ULA
END BEHAVIORAL;

