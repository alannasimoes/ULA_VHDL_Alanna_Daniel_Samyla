--------------------------------------------------------------------------------
-- COMPANY: 
-- ENGINEER:
--
-- CREATE DATE:   00:33:46 06/18/2024
-- DESIGN NAME:   
-- MODULE NAME:   C:/USERS/DANIEL/DESKTOP/SD/ULA_FINAL/TB_ULA.VHD
-- PROJECT NAME:  ULA_FINAL
-- TARGET DEVICE:  
-- TOOL VERSIONS:  
-- DESCRIPTION:   
-- 
-- VHDL TEST BENCH CREATED BY ISE FOR MODULE: ULA
-- 
-- DEPENDENCIES:
-- 
-- REVISION:
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS:
--
-- NOTES: 
-- THIS TESTBENCH HAS BEEN AUTOMATICALLY GENERATED USING TYPES STD_LOGIC AND
-- STD_LOGIC_VECTOR FOR THE PORTS OF THE UNIT UNDER TEST.  XILINX RECOMMENDS
-- THAT THESE TYPES ALWAYS BE USED FOR THE TOP-LEVEL I/O OF A DESIGN IN ORDER
-- TO GUARANTEE THAT THE TESTBENCH WILL BIND CORRECTLY TO THE POST-IMPLEMENTATION 
-- SIMULATION MODEL.
--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 
-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;
 
ENTITY TB_ULA IS
END TB_ULA;
 
ARCHITECTURE BEHAVIOR OF TB_ULA IS 
 
    -- COMPONENT DECLARATION FOR THE UNIT UNDER TEST (UUT)
 
    COMPONENT ULA
    PORT(
         A_ULA : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         B_ULA : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         SEL_ULA : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
         RESULTADO_ULA : OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
         FLAG_CARRY_OUT_ULA : OUT  STD_LOGIC;
         FLAG_RESULTADO_NULO_ULA : OUT  STD_LOGIC;
         FLAG_OVERFLOW_ULA : OUT  STD_LOGIC;
			FLAG_RESULTADO_NEGATIVO_ULA : OUT  STD_LOGIC
        );
    END COMPONENT;
    

   --INPUTS
   SIGNAL A_ULA : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
   SIGNAL B_ULA : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
   SIGNAL SEL_ULA : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');

 	--OUTPUTS
   SIGNAL RESULTADO_ULA : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL FLAG_CARRY_OUT_ULA : STD_LOGIC;
   SIGNAL FLAG_RESULTADO_NULO_ULA : STD_LOGIC;
   SIGNAL FLAG_OVERFLOW_ULA : STD_LOGIC;
	SIGNAL FLAG_RESULTADO_NEGATIVO_ULA : STD_LOGIC;
 
BEGIN
 
	-- INSTANTIATE THE UNIT UNDER TEST (UUT)
   UUT: ULA PORT MAP (
          A_ULA => A_ULA,
          B_ULA => B_ULA,
          SEL_ULA => SEL_ULA,
          RESULTADO_ULA => RESULTADO_ULA,
          FLAG_CARRY_OUT_ULA => FLAG_CARRY_OUT_ULA,
          FLAG_RESULTADO_NULO_ULA => FLAG_RESULTADO_NULO_ULA,
          FLAG_OVERFLOW_ULA => FLAG_OVERFLOW_ULA,
			 FLAG_RESULTADO_NEGATIVO_ULA => FLAG_RESULTADO_NEGATIVO_ULA
        );

 
-- STIMULUS PROCESS
   STIM_PROC: PROCESS
   BEGIN
		--- TESTE DE AND
		A_ULA <= "0001";
		B_ULA <= "0001";
		SEL_ULA <= "000";
		WAIT FOR 100 NS;
		--- TESTE DE OR
		A_ULA <= "0000";
		B_ULA <= "0001";
		SEL_ULA <= "001";
		WAIT FOR 100 NS;
		--- TESTE DE NOT
		A_ULA <= "0000";
		B_ULA <= "0001";
		SEL_ULA <= "010";
		WAIT FOR 100 NS;
		--- TESTE DE XOR
		A_ULA <= "0000";
		B_ULA <= "0000";
		SEL_ULA <= "011";
		WAIT FOR 100 NS;
		--- TESTE DE SOMA
		A_ULA <= "1111";
		B_ULA <= "0001";
		SEL_ULA <= "100";
		WAIT FOR 100 NS;
		--- TESTE DE SUBTRACAO
		A_ULA <= "0010";
		B_ULA <= "0100";
		SEL_ULA <= "101";
		WAIT FOR 100 NS;
		--- TESTE DE COMPARACAO
		A_ULA <= "0100";
		B_ULA <= "0010";
		SEL_ULA <= "110";
		--- TESTE DE DESLOCAMENTO
		A_ULA <= "0100";
		SEL_ULA <= "111";
		WAIT FOR 100 NS;
      WAIT;
   END PROCESS;


END;
